module server_time

fn test_get() {
  println(get('testnet.binance.vision')!)
}
